package Synchronous_FIFO_package;

`include "Synchronous_FIFO_transaction.sv"
`include "Synchronous_FIFO_generator.sv"
`include "Synchronous_FIFO_driver.sv"
`include "Synchronous_FIFO_monitor.sv"
`include "Synchronous_FIFO_scoreboard.sv"
`include "Synchronous_FIFO_env.sv"

endpackage
